VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DIGITALTBD
  CLASS BLOCK ;
  FOREIGN DIGITALTBD ;
  ORIGIN 0.000 0.000 ;
  
  # Reduced from `caravel_user` by (10x10)um (5um per side)
  SIZE 2910.000 BY 3510.000 ;

  PIN VCCD1
    PORT
      LAYER met3 ;
        RECT 2833.630 3193.920 2924.000 3217.920 ;
    END
  END VCCD1
  PIN VDDA1
    PORT
      LAYER met3 ;
        RECT 2811.595 2747.810 2924.000 2771.810 ;
    END
  END VDDA1
  PIN VSSA1
    PORT
      LAYER met3 ;
        RECT 2547.970 3182.805 2571.970 3416.680 ;
    END
  END VSSA1
  PIN VSSD1
    PORT
      LAYER met3 ;
        RECT 82.105 952.150 2863.025 976.150 ;
    END
  END VSSD1
  PIN gpio_analog[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1341.150 2924.000 1341.710 ;
    END
  END gpio_analog[0]
  PIN gpio_analog[10]
    PORT
      LAYER met3 ;
        RECT -14.000 1904.320 -7.600 1904.880 ;
    END
  END gpio_analog[10]
  PIN gpio_analog[11]
    PORT
      LAYER met3 ;
        RECT -14.000 1688.210 -7.600 1688.770 ;
    END
  END gpio_analog[11]
  PIN gpio_analog[12]
    PORT
      LAYER met3 ;
        RECT -14.000 1472.100 -7.600 1472.660 ;
    END
  END gpio_analog[12]
  PIN gpio_analog[13]
    PORT
      LAYER met3 ;
        RECT -14.000 1256.990 -7.600 1257.550 ;
    END
  END gpio_analog[13]
  PIN gpio_analog[14]
    PORT
      LAYER met3 ;
        RECT -14.000 618.880 -7.600 619.440 ;
    END
  END gpio_analog[14]
  PIN gpio_analog[15]
    PORT
      LAYER met3 ;
        RECT -14.000 402.770 -7.600 403.330 ;
    END
  END gpio_analog[15]
  PIN gpio_analog[16]
    PORT
      LAYER met3 ;
        RECT -14.000 186.660 -7.600 187.220 ;
    END
  END gpio_analog[16]
  PIN gpio_analog[17]
    PORT
      LAYER met3 ;
        RECT -14.000 79.550 -7.600 80.110 ;
    END
  END gpio_analog[17]
  PIN gpio_analog[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1563.260 2924.000 1563.820 ;
    END
  END gpio_analog[1]
  PIN gpio_analog[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1789.370 2924.000 1789.930 ;
    END
  END gpio_analog[2]
  PIN gpio_analog[3]
    PORT
      LAYER met3 ;
        RECT 2667.485 2021.480 2924.000 2022.040 ;
    END
  END gpio_analog[3]
  PIN gpio_analog[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2243.590 2924.000 2244.150 ;
    END
  END gpio_analog[4]
  PIN gpio_analog[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2465.700 2924.000 2466.260 ;
    END
  END gpio_analog[5]
  PIN gpio_analog[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2912.810 2924.000 2913.370 ;
    END
  END gpio_analog[6]
  PIN gpio_analog[7]
    PORT
      LAYER met3 ;
        RECT -14.000 2552.650 1690.360 2553.210 ;
    END
  END gpio_analog[7]
  PIN gpio_analog[8]
    PORT
      LAYER met3 ;
        RECT -14.000 2336.540 -7.600 2337.100 ;
    END
  END gpio_analog[8]
  PIN gpio_analog[9]
    PORT
      LAYER met3 ;
        RECT -14.000 2120.430 -7.600 2120.990 ;
    END
  END gpio_analog[9]
  PIN gpio_noesd[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1347.060 2924.000 1347.620 ;
    END
  END gpio_noesd[0]
  PIN gpio_noesd[10]
    PORT
      LAYER met3 ;
        RECT -14.000 1898.410 -7.600 1898.970 ;
    END
  END gpio_noesd[10]
  PIN gpio_noesd[11]
    PORT
      LAYER met3 ;
        RECT -14.000 1682.300 -7.600 1682.860 ;
    END
  END gpio_noesd[11]
  PIN gpio_noesd[12]
    PORT
      LAYER met3 ;
        RECT -14.000 1466.190 -7.600 1466.750 ;
    END
  END gpio_noesd[12]
  PIN gpio_noesd[13]
    PORT
      LAYER met3 ;
        RECT -14.000 1251.080 -7.600 1251.640 ;
    END
  END gpio_noesd[13]
  PIN gpio_noesd[14]
    PORT
      LAYER met3 ;
        RECT -14.000 612.970 -7.600 613.530 ;
    END
  END gpio_noesd[14]
  PIN gpio_noesd[15]
    PORT
      LAYER met3 ;
        RECT -14.000 396.860 -7.600 397.420 ;
    END
  END gpio_noesd[15]
  PIN gpio_noesd[16]
    PORT
      LAYER met3 ;
        RECT -14.000 180.750 -7.600 181.310 ;
    END
  END gpio_noesd[16]
  PIN gpio_noesd[17]
    PORT
      LAYER met3 ;
        RECT -14.000 73.640 -7.600 74.200 ;
    END
  END gpio_noesd[17]
  PIN gpio_noesd[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1569.170 2924.000 1569.730 ;
    END
  END gpio_noesd[1]
  PIN gpio_noesd[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1795.280 2924.000 1795.840 ;
    END
  END gpio_noesd[2]
  PIN gpio_noesd[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 2027.390 2924.000 2027.950 ;
    END
  END gpio_noesd[3]
  PIN gpio_noesd[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2249.500 2924.000 2250.060 ;
    END
  END gpio_noesd[4]
  PIN gpio_noesd[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2471.610 2924.000 2472.170 ;
    END
  END gpio_noesd[5]
  PIN gpio_noesd[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2918.720 2924.000 2919.280 ;
    END
  END gpio_noesd[6]
  PIN gpio_noesd[7]
    PORT
      LAYER met3 ;
        RECT -14.000 2546.740 -7.600 2547.300 ;
    END
  END gpio_noesd[7]
  PIN gpio_noesd[8]
    PORT
      LAYER met3 ;
        RECT -14.000 2330.630 -7.600 2331.190 ;
    END
  END gpio_noesd[8]
  PIN gpio_noesd[9]
    PORT
      LAYER met3 ;
        RECT -14.000 2114.520 -7.600 2115.080 ;
    END
  END gpio_noesd[9]
  PIN io_analog[0]
    PORT
      LAYER met3 ;
        RECT 2911.500 3384.920 2924.000 3409.920 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    PORT
      LAYER met3 ;
        RECT -14.000 3396.210 -1.500 3421.210 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    PORT
      LAYER met3 ;
        RECT 2827.970 3501.500 2852.970 3514.000 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    PORT
      LAYER met3 ;
        RECT 2321.970 3501.500 2346.970 3514.000 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    PORT
      LAYER met3 ;
        RECT 2061.970 3501.500 2086.970 3514.000 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    PORT
      LAYER met3 ;
        RECT 1641.470 3237.450 1666.470 3514.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1589.970 3237.450 1614.970 3514.000 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    PORT
      LAYER met3 ;
        RECT 1132.970 3501.500 1157.970 3514.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1081.470 3501.500 1106.470 3514.000 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    PORT
      LAYER met3 ;
        RECT 874.470 3501.500 899.470 3514.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 822.970 3501.500 847.970 3514.000 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    PORT
      LAYER met3 ;
        RECT 595.970 3501.500 620.970 3514.000 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    PORT
      LAYER met3 ;
        RECT 335.970 3501.500 360.970 3514.000 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    PORT
      LAYER met3 ;
        RECT 75.970 3501.500 100.970 3514.000 ;
    END
  END io_analog[9]
  PIN io_clamp_high[0]
    PORT
      LAYER met3 ;
        RECT 1628.970 3450.460 1639.970 3514.000 ;
    END
  END io_clamp_high[0]
  PIN io_clamp_high[1]
    PORT
      LAYER met3 ;
        RECT 1120.470 3443.050 1131.470 3514.000 ;
    END
  END io_clamp_high[1]
  PIN io_clamp_high[2]
    PORT
      LAYER met3 ;
        RECT 861.970 3442.885 872.970 3514.000 ;
    END
  END io_clamp_high[2]
  PIN io_clamp_low[0]
    PORT
      LAYER met3 ;
        RECT 1616.470 3442.965 1627.470 3514.000 ;
    END
  END io_clamp_low[0]
  PIN io_clamp_low[1]
    PORT
      LAYER met3 ;
        RECT 1107.970 3443.050 1118.970 3514.000 ;
    END
  END io_clamp_low[1]
  PIN io_clamp_low[2]
    PORT
      LAYER met3 ;
        RECT 849.470 3442.885 860.470 3514.000 ;
    END
  END io_clamp_low[2]
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 8.630 2924.000 9.190 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2039.210 2924.000 2039.770 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2261.320 2924.000 2261.880 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2483.430 2924.000 2483.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2930.540 2924.000 2931.100 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met3 ;
        RECT -14.000 2534.920 -7.600 2535.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met3 ;
        RECT -14.000 2318.810 -7.600 2319.370 ;
    END
  END io_in[15]
  PIN io_in[16]
    PORT
      LAYER met3 ;
        RECT -14.000 2102.700 -7.600 2103.260 ;
    END
  END io_in[16]
  PIN io_in[17]
    PORT
      LAYER met3 ;
        RECT -14.000 1886.590 -7.600 1887.150 ;
    END
  END io_in[17]
  PIN io_in[18]
    PORT
      LAYER met3 ;
        RECT -14.000 1670.480 -7.600 1671.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    PORT
      LAYER met3 ;
        RECT -14.000 1454.370 -7.600 1454.930 ;
    END
  END io_in[19]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 32.270 2924.000 32.830 ;
    END
  END io_in[1]
  PIN io_in[20]
    PORT
      LAYER met3 ;
        RECT -14.000 1239.260 -7.600 1239.820 ;
    END
  END io_in[20]
  PIN io_in[21]
    PORT
      LAYER met3 ;
        RECT -14.000 601.150 -7.600 601.710 ;
    END
  END io_in[21]
  PIN io_in[22]
    PORT
      LAYER met3 ;
        RECT -14.000 385.040 -7.600 385.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    PORT
      LAYER met3 ;
        RECT -14.000 168.930 -7.600 169.490 ;
    END
  END io_in[23]
  PIN io_in[24]
    PORT
      LAYER met3 ;
        RECT -14.000 61.820 -7.600 62.380 ;
    END
  END io_in[24]
  PIN io_in[25]
    PORT
      LAYER met3 ;
        RECT -14.000 38.180 -7.600 38.740 ;
    END
  END io_in[25]
  PIN io_in[26]
    PORT
      LAYER met3 ;
        RECT -14.000 14.540 -7.600 15.100 ;
    END
  END io_in[26]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 55.910 2924.000 56.470 ;
    END
  END io_in[2]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 79.550 2924.000 80.110 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 103.190 2924.000 103.750 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 235.480 2924.000 236.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 458.770 2924.000 459.330 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1358.880 2924.000 1359.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1580.990 2924.000 1581.550 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1807.100 2924.000 1807.660 ;
    END
  END io_in[9]
  PIN io_in_3v3[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 2.720 2924.000 3.280 ;
    END
  END io_in_3v3[0]
  PIN io_in_3v3[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2033.300 2924.000 2033.860 ;
    END
  END io_in_3v3[10]
  PIN io_in_3v3[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2255.410 2924.000 2255.970 ;
    END
  END io_in_3v3[11]
  PIN io_in_3v3[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2477.520 2924.000 2478.080 ;
    END
  END io_in_3v3[12]
  PIN io_in_3v3[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2924.630 2924.000 2925.190 ;
    END
  END io_in_3v3[13]
  PIN io_in_3v3[14]
    PORT
      LAYER met3 ;
        RECT -14.000 2540.830 -7.600 2541.390 ;
    END
  END io_in_3v3[14]
  PIN io_in_3v3[15]
    PORT
      LAYER met3 ;
        RECT -14.000 2324.720 -7.600 2325.280 ;
    END
  END io_in_3v3[15]
  PIN io_in_3v3[16]
    PORT
      LAYER met3 ;
        RECT -14.000 2108.610 -7.600 2109.170 ;
    END
  END io_in_3v3[16]
  PIN io_in_3v3[17]
    PORT
      LAYER met3 ;
        RECT -14.000 1892.500 -7.600 1893.060 ;
    END
  END io_in_3v3[17]
  PIN io_in_3v3[18]
    PORT
      LAYER met3 ;
        RECT -14.000 1676.390 -7.600 1676.950 ;
    END
  END io_in_3v3[18]
  PIN io_in_3v3[19]
    PORT
      LAYER met3 ;
        RECT -14.000 1460.280 -7.600 1460.840 ;
    END
  END io_in_3v3[19]
  PIN io_in_3v3[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 26.360 2924.000 26.920 ;
    END
  END io_in_3v3[1]
  PIN io_in_3v3[20]
    PORT
      LAYER met3 ;
        RECT -14.000 1245.170 -7.600 1245.730 ;
    END
  END io_in_3v3[20]
  PIN io_in_3v3[21]
    PORT
      LAYER met3 ;
        RECT -14.000 607.060 -7.600 607.620 ;
    END
  END io_in_3v3[21]
  PIN io_in_3v3[22]
    PORT
      LAYER met3 ;
        RECT -14.000 390.950 -7.600 391.510 ;
    END
  END io_in_3v3[22]
  PIN io_in_3v3[23]
    PORT
      LAYER met3 ;
        RECT -14.000 174.840 -7.600 175.400 ;
    END
  END io_in_3v3[23]
  PIN io_in_3v3[24]
    PORT
      LAYER met3 ;
        RECT -14.000 67.730 -7.600 68.290 ;
    END
  END io_in_3v3[24]
  PIN io_in_3v3[25]
    PORT
      LAYER met3 ;
        RECT -14.000 44.090 -7.600 44.650 ;
    END
  END io_in_3v3[25]
  PIN io_in_3v3[26]
    PORT
      LAYER met3 ;
        RECT -14.000 20.450 -7.600 21.010 ;
    END
  END io_in_3v3[26]
  PIN io_in_3v3[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 50.000 2924.000 50.560 ;
    END
  END io_in_3v3[2]
  PIN io_in_3v3[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 73.640 2924.000 74.200 ;
    END
  END io_in_3v3[3]
  PIN io_in_3v3[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 97.280 2924.000 97.840 ;
    END
  END io_in_3v3[4]
  PIN io_in_3v3[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 229.570 2924.000 230.130 ;
    END
  END io_in_3v3[5]
  PIN io_in_3v3[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 452.860 2924.000 453.420 ;
    END
  END io_in_3v3[6]
  PIN io_in_3v3[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1352.970 2924.000 1353.530 ;
    END
  END io_in_3v3[7]
  PIN io_in_3v3[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1575.080 2924.000 1575.640 ;
    END
  END io_in_3v3[8]
  PIN io_in_3v3[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1801.190 2924.000 1801.750 ;
    END
  END io_in_3v3[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 20.450 2924.000 21.010 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2051.030 2924.000 2051.590 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met3 ;
        RECT 2898.095 2273.140 2924.000 2273.700 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met3 ;
        RECT 2898.095 2495.250 2924.000 2495.810 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2942.360 2924.000 2942.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT -14.000 2523.100 -7.600 2523.660 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met3 ;
        RECT -14.000 2306.990 59.485 2307.550 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    PORT
      LAYER met3 ;
        RECT -14.000 2090.880 59.555 2091.440 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    PORT
      LAYER met3 ;
        RECT -14.000 1874.770 -7.600 1875.330 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    PORT
      LAYER met3 ;
        RECT -14.000 1658.660 -7.600 1659.220 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    PORT
      LAYER met3 ;
        RECT -14.000 1442.550 -7.600 1443.110 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 44.090 2924.000 44.650 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    PORT
      LAYER met3 ;
        RECT -14.000 1227.440 -7.600 1228.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    PORT
      LAYER met3 ;
        RECT -14.000 589.330 -7.600 589.890 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    PORT
      LAYER met3 ;
        RECT -14.000 373.220 -7.600 373.780 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    PORT
      LAYER met3 ;
        RECT -14.000 157.110 -7.600 157.670 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    PORT
      LAYER met3 ;
        RECT -14.000 50.000 -7.600 50.560 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    PORT
      LAYER met3 ;
        RECT -14.000 26.360 -7.600 26.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    PORT
      LAYER met3 ;
        RECT -14.000 2.720 -7.600 3.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 67.730 2924.000 68.290 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 91.370 2924.000 91.930 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 115.010 2924.000 115.570 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 247.300 2924.000 247.860 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 470.590 2924.000 471.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1370.700 2924.000 1371.260 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1592.810 2924.000 1593.370 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1818.920 2924.000 1819.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 14.540 2924.000 15.100 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2045.120 2924.000 2045.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 2686.880 2267.230 2924.000 2267.790 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT 2697.470 2489.340 2924.000 2489.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2936.450 2924.000 2937.010 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met3 ;
        RECT -14.000 2529.010 -7.600 2529.570 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met3 ;
        RECT -14.000 2312.900 1695.395 2313.460 ;
    END
  END io_out[15]
  PIN io_out[16]
    PORT
      LAYER met3 ;
        RECT -14.000 2096.790 1699.250 2097.350 ;
    END
  END io_out[16]
  PIN io_out[17]
    PORT
      LAYER met3 ;
        RECT -14.000 1880.680 -7.600 1881.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    PORT
      LAYER met3 ;
        RECT -14.000 1664.570 -7.600 1665.130 ;
    END
  END io_out[18]
  PIN io_out[19]
    PORT
      LAYER met3 ;
        RECT -14.000 1448.460 -7.600 1449.020 ;
    END
  END io_out[19]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 38.180 2924.000 38.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    PORT
      LAYER met3 ;
        RECT -14.000 1233.350 -7.600 1233.910 ;
    END
  END io_out[20]
  PIN io_out[21]
    PORT
      LAYER met3 ;
        RECT -14.000 595.240 -7.600 595.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    PORT
      LAYER met3 ;
        RECT -14.000 379.130 -7.600 379.690 ;
    END
  END io_out[22]
  PIN io_out[23]
    PORT
      LAYER met3 ;
        RECT -14.000 163.020 -7.600 163.580 ;
    END
  END io_out[23]
  PIN io_out[24]
    PORT
      LAYER met3 ;
        RECT -14.000 55.910 -7.600 56.470 ;
    END
  END io_out[24]
  PIN io_out[25]
    PORT
      LAYER met3 ;
        RECT -14.000 32.270 -7.600 32.830 ;
    END
  END io_out[25]
  PIN io_out[26]
    PORT
      LAYER met3 ;
        RECT -14.000 8.630 -7.600 9.190 ;
    END
  END io_out[26]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 61.820 2924.000 62.380 ;
    END
  END io_out[2]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 85.460 2924.000 86.020 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 109.100 2924.000 109.660 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 241.390 2924.000 241.950 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 464.680 2924.000 465.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1364.790 2924.000 1365.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1586.900 2924.000 1587.460 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1813.010 2924.000 1813.570 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 624.080 -4.000 624.640 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met2 ;
        RECT 2397.080 -4.000 2397.640 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met2 ;
        RECT 2414.810 -4.000 2415.370 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 2432.540 -4.000 2433.100 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met2 ;
        RECT 2450.270 -4.000 2450.830 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met2 ;
        RECT 2468.000 -4.000 2468.560 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 2485.730 -4.000 2486.290 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 2503.460 -4.000 2504.020 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met2 ;
        RECT 2521.190 -4.000 2521.750 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met2 ;
        RECT 2538.920 -4.000 2539.480 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met2 ;
        RECT 2556.650 -4.000 2557.210 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met2 ;
        RECT 801.380 -4.000 801.940 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met2 ;
        RECT 2574.380 -4.000 2574.940 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met2 ;
        RECT 2592.110 -4.000 2592.670 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met2 ;
        RECT 2609.840 -4.000 2610.400 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met2 ;
        RECT 2627.570 -4.000 2628.130 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met2 ;
        RECT 2645.300 -4.000 2645.860 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 2663.030 -4.000 2663.590 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 2680.760 -4.000 2681.320 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met2 ;
        RECT 2698.490 -4.000 2699.050 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met2 ;
        RECT 2716.220 -4.000 2716.780 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met2 ;
        RECT 2733.950 -4.000 2734.510 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 819.110 -4.000 819.670 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met2 ;
        RECT 2751.680 -4.000 2752.240 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 2769.410 -4.000 2769.970 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 2787.140 -4.000 2787.700 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met2 ;
        RECT 2804.870 -4.000 2805.430 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 2822.600 -4.000 2823.160 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 2840.330 -4.000 2840.890 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met2 ;
        RECT 2858.060 -4.000 2858.620 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2875.790 -4.000 2876.350 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met2 ;
        RECT 836.840 -4.000 837.400 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met2 ;
        RECT 854.570 -4.000 855.130 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met2 ;
        RECT 872.300 -4.000 872.860 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met2 ;
        RECT 890.030 -4.000 890.590 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met2 ;
        RECT 907.760 -4.000 908.320 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met2 ;
        RECT 925.490 -4.000 926.050 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met2 ;
        RECT 943.220 -4.000 943.780 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 960.950 -4.000 961.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 641.810 -4.000 642.370 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met2 ;
        RECT 978.680 -4.000 979.240 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 996.410 -4.000 996.970 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 1014.140 -4.000 1014.700 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met2 ;
        RECT 1031.870 -4.000 1032.430 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met2 ;
        RECT 1049.600 -4.000 1050.160 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 1067.330 -4.000 1067.890 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 1085.060 -4.000 1085.620 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 1102.790 -4.000 1103.350 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met2 ;
        RECT 1120.520 -4.000 1121.080 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met2 ;
        RECT 1138.250 -4.000 1138.810 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 659.540 -4.000 660.100 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met2 ;
        RECT 1155.980 -4.000 1156.540 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met2 ;
        RECT 1173.710 -4.000 1174.270 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 1191.440 -4.000 1192.000 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met2 ;
        RECT 1209.170 -4.000 1209.730 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met2 ;
        RECT 1226.900 -4.000 1227.460 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met2 ;
        RECT 1244.630 -4.000 1245.190 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 1262.360 -4.000 1262.920 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 1280.090 -4.000 1280.650 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 1297.820 -4.000 1298.380 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 1315.550 -4.000 1316.110 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met2 ;
        RECT 677.270 -4.000 677.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 1333.280 -4.000 1333.840 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met2 ;
        RECT 1351.010 -4.000 1351.570 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met2 ;
        RECT 1368.740 -4.000 1369.300 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met2 ;
        RECT 1386.470 -4.000 1387.030 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met2 ;
        RECT 1404.200 -4.000 1404.760 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 1421.930 -4.000 1422.490 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 1439.660 -4.000 1440.220 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met2 ;
        RECT 1457.390 -4.000 1457.950 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met2 ;
        RECT 1475.120 -4.000 1475.680 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met2 ;
        RECT 1492.850 -4.000 1493.410 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 695.000 -4.000 695.560 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 1510.580 -4.000 1511.140 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met2 ;
        RECT 1528.310 -4.000 1528.870 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met2 ;
        RECT 1546.040 -4.000 1546.600 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 1563.770 -4.000 1564.330 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 1581.500 -4.000 1582.060 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met2 ;
        RECT 1599.230 -4.000 1599.790 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met2 ;
        RECT 1616.960 -4.000 1617.520 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met2 ;
        RECT 1634.690 -4.000 1635.250 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 1652.420 -4.000 1652.980 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met2 ;
        RECT 1670.150 -4.000 1670.710 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met2 ;
        RECT 712.730 -4.000 713.290 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 1687.880 -4.000 1688.440 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 1705.610 -4.000 1706.170 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met2 ;
        RECT 1723.340 -4.000 1723.900 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met2 ;
        RECT 1741.070 -4.000 1741.630 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met2 ;
        RECT 1758.800 -4.000 1759.360 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met2 ;
        RECT 1776.530 -4.000 1777.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met2 ;
        RECT 1794.260 -4.000 1794.820 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 1811.990 -4.000 1812.550 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met2 ;
        RECT 1829.720 -4.000 1830.280 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met2 ;
        RECT 1847.450 -4.000 1848.010 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met2 ;
        RECT 730.460 -4.000 731.020 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met2 ;
        RECT 1865.180 -4.000 1865.740 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met2 ;
        RECT 1882.910 -4.000 1883.470 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 1900.640 -4.000 1901.200 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met2 ;
        RECT 1918.370 -4.000 1918.930 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met2 ;
        RECT 1936.100 -4.000 1936.660 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 1953.830 -4.000 1954.390 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met2 ;
        RECT 1971.560 -4.000 1972.120 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 1989.290 -4.000 1989.850 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 2007.020 -4.000 2007.580 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met2 ;
        RECT 2024.750 -4.000 2025.310 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 748.190 -4.000 748.750 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met2 ;
        RECT 2042.480 -4.000 2043.040 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 2060.210 -4.000 2060.770 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 2077.940 -4.000 2078.500 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met2 ;
        RECT 2095.670 -4.000 2096.230 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met2 ;
        RECT 2113.400 -4.000 2113.960 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met2 ;
        RECT 2131.130 -4.000 2131.690 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met2 ;
        RECT 2148.860 -4.000 2149.420 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 2166.590 -4.000 2167.150 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met2 ;
        RECT 2184.320 -4.000 2184.880 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 2202.050 -4.000 2202.610 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 765.920 -4.000 766.480 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met2 ;
        RECT 2219.780 -4.000 2220.340 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met2 ;
        RECT 2237.510 -4.000 2238.070 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met2 ;
        RECT 2255.240 -4.000 2255.800 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met2 ;
        RECT 2272.970 -4.000 2273.530 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met2 ;
        RECT 2290.700 -4.000 2291.260 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met2 ;
        RECT 2308.430 -4.000 2308.990 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met2 ;
        RECT 2326.160 -4.000 2326.720 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met2 ;
        RECT 2343.890 -4.000 2344.450 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 2361.620 -4.000 2362.180 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met2 ;
        RECT 2379.350 -4.000 2379.910 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 783.650 -4.000 784.210 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met2 ;
        RECT 629.990 -4.000 630.550 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 2402.990 -4.000 2403.550 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 2420.720 -4.000 2421.280 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 2438.450 -4.000 2439.010 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met2 ;
        RECT 2456.180 -4.000 2456.740 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 2473.910 -4.000 2474.470 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met2 ;
        RECT 2491.640 -4.000 2492.200 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 2509.370 -4.000 2509.930 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met2 ;
        RECT 2527.100 -4.000 2527.660 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met2 ;
        RECT 2544.830 -4.000 2545.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 2562.560 -4.000 2563.120 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met2 ;
        RECT 807.290 -4.000 807.850 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met2 ;
        RECT 2580.290 -4.000 2580.850 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met2 ;
        RECT 2598.020 -4.000 2598.580 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met2 ;
        RECT 2615.750 -4.000 2616.310 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 2633.480 -4.000 2634.040 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 2651.210 -4.000 2651.770 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 2668.940 -4.000 2669.500 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 2686.670 -4.000 2687.230 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met2 ;
        RECT 2704.400 -4.000 2704.960 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met2 ;
        RECT 2722.130 -4.000 2722.690 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met2 ;
        RECT 2739.860 -4.000 2740.420 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 825.020 -4.000 825.580 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 2757.590 -4.000 2758.150 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 2775.320 -4.000 2775.880 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 2793.050 -4.000 2793.610 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met2 ;
        RECT 2810.780 -4.000 2811.340 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met2 ;
        RECT 2828.510 -4.000 2829.070 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met2 ;
        RECT 2846.240 -4.000 2846.800 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met2 ;
        RECT 2863.970 -4.000 2864.530 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met2 ;
        RECT 2881.700 -4.000 2882.260 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 842.750 -4.000 843.310 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met2 ;
        RECT 860.480 -4.000 861.040 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met2 ;
        RECT 878.210 -4.000 878.770 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met2 ;
        RECT 895.940 -4.000 896.500 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 913.670 -4.000 914.230 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met2 ;
        RECT 931.400 -4.000 931.960 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 949.130 -4.000 949.690 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 966.860 -4.000 967.420 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met2 ;
        RECT 647.720 -4.000 648.280 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met2 ;
        RECT 984.590 -4.000 985.150 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met2 ;
        RECT 1002.320 -4.000 1002.880 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met2 ;
        RECT 1020.050 -4.000 1020.610 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met2 ;
        RECT 1037.780 -4.000 1038.340 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met2 ;
        RECT 1055.510 -4.000 1056.070 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 1073.240 -4.000 1073.800 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met2 ;
        RECT 1090.970 -4.000 1091.530 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met2 ;
        RECT 1108.700 -4.000 1109.260 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 1126.430 -4.000 1126.990 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 1144.160 -4.000 1144.720 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 665.450 -4.000 666.010 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 1161.890 -4.000 1162.450 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met2 ;
        RECT 1179.620 -4.000 1180.180 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met2 ;
        RECT 1197.350 -4.000 1197.910 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met2 ;
        RECT 1215.080 -4.000 1215.640 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 1232.810 -4.000 1233.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met2 ;
        RECT 1250.540 -4.000 1251.100 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 1268.270 -4.000 1268.830 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met2 ;
        RECT 1286.000 -4.000 1286.560 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met2 ;
        RECT 1303.730 -4.000 1304.290 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met2 ;
        RECT 1321.460 -4.000 1322.020 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met2 ;
        RECT 683.180 -4.000 683.740 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met2 ;
        RECT 1339.190 -4.000 1339.750 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 1356.920 -4.000 1357.480 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 1374.650 -4.000 1375.210 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met2 ;
        RECT 1392.380 -4.000 1392.940 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 1410.110 -4.000 1410.670 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 1427.840 -4.000 1428.400 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 1445.570 -4.000 1446.130 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met2 ;
        RECT 1463.300 -4.000 1463.860 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 1481.030 -4.000 1481.590 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 1498.760 -4.000 1499.320 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 700.910 -4.000 701.470 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met2 ;
        RECT 1516.490 -4.000 1517.050 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 1534.220 -4.000 1534.780 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met2 ;
        RECT 1551.950 -4.000 1552.510 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 1569.680 -4.000 1570.240 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 1587.410 -4.000 1587.970 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met2 ;
        RECT 1605.140 -4.000 1605.700 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 1622.870 -4.000 1623.430 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 1640.600 -4.000 1641.160 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met2 ;
        RECT 1658.330 -4.000 1658.890 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met2 ;
        RECT 1676.060 -4.000 1676.620 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 718.640 -4.000 719.200 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met2 ;
        RECT 1693.790 -4.000 1694.350 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met2 ;
        RECT 1711.520 -4.000 1712.080 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1729.250 -4.000 1729.810 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 1746.980 -4.000 1747.540 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met2 ;
        RECT 1764.710 -4.000 1765.270 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 1782.440 -4.000 1783.000 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met2 ;
        RECT 1800.170 -4.000 1800.730 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met2 ;
        RECT 1817.900 -4.000 1818.460 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met2 ;
        RECT 1835.630 -4.000 1836.190 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met2 ;
        RECT 1853.360 -4.000 1853.920 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 736.370 -4.000 736.930 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 1871.090 -4.000 1871.650 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met2 ;
        RECT 1888.820 -4.000 1889.380 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 1906.550 -4.000 1907.110 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1924.280 -4.000 1924.840 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 1942.010 -4.000 1942.570 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 1959.740 -4.000 1960.300 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met2 ;
        RECT 1977.470 -4.000 1978.030 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met2 ;
        RECT 1995.200 -4.000 1995.760 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 2012.930 -4.000 2013.490 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met2 ;
        RECT 2030.660 -4.000 2031.220 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met2 ;
        RECT 754.100 -4.000 754.660 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met2 ;
        RECT 2048.390 -4.000 2048.950 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met2 ;
        RECT 2066.120 -4.000 2066.680 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 2083.850 -4.000 2084.410 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met2 ;
        RECT 2101.580 -4.000 2102.140 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 2119.310 -4.000 2119.870 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 2137.040 -4.000 2137.600 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 2154.770 -4.000 2155.330 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 2172.500 -4.000 2173.060 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met2 ;
        RECT 2190.230 -4.000 2190.790 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met2 ;
        RECT 2207.960 -4.000 2208.520 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met2 ;
        RECT 771.830 -4.000 772.390 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 2225.690 -4.000 2226.250 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 2243.420 -4.000 2243.980 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 2261.150 -4.000 2261.710 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 2278.880 -4.000 2279.440 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 2296.610 -4.000 2297.170 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met2 ;
        RECT 2314.340 -4.000 2314.900 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 2332.070 -4.000 2332.630 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 2349.800 -4.000 2350.360 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 2367.530 -4.000 2368.090 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 2385.260 -4.000 2385.820 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met2 ;
        RECT 789.560 -4.000 790.120 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 635.900 -4.000 636.460 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met2 ;
        RECT 2408.900 -4.000 2409.460 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met2 ;
        RECT 2426.630 -4.000 2427.190 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 2444.360 -4.000 2444.920 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 2462.090 -4.000 2462.650 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 2479.820 -4.000 2480.380 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met2 ;
        RECT 2497.550 -4.000 2498.110 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 2515.280 -4.000 2515.840 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 2533.010 -4.000 2533.570 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met2 ;
        RECT 2550.740 -4.000 2551.300 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 2568.470 -4.000 2569.030 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 813.200 -4.000 813.760 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 2586.200 -4.000 2586.760 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 2603.930 -4.000 2604.490 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met2 ;
        RECT 2621.660 -4.000 2622.220 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 2639.390 -4.000 2639.950 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met2 ;
        RECT 2657.120 -4.000 2657.680 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 2674.850 -4.000 2675.410 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met2 ;
        RECT 2692.580 -4.000 2693.140 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 2710.310 -4.000 2710.870 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 2728.040 -4.000 2728.600 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met2 ;
        RECT 2745.770 -4.000 2746.330 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 830.930 -4.000 831.490 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 2763.500 -4.000 2764.060 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met2 ;
        RECT 2781.230 -4.000 2781.790 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met2 ;
        RECT 2798.960 -4.000 2799.520 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 2816.690 -4.000 2817.250 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 2834.420 -4.000 2834.980 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 2852.150 -4.000 2852.710 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 2869.880 -4.000 2870.440 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met2 ;
        RECT 2887.610 -4.000 2888.170 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met2 ;
        RECT 848.660 -4.000 849.220 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met2 ;
        RECT 866.390 -4.000 866.950 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met2 ;
        RECT 884.120 -4.000 884.680 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met2 ;
        RECT 901.850 -4.000 902.410 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met2 ;
        RECT 919.580 -4.000 920.140 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 937.310 -4.000 937.870 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met2 ;
        RECT 955.040 -4.000 955.600 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met2 ;
        RECT 972.770 -4.000 973.330 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 653.630 -4.000 654.190 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met2 ;
        RECT 990.500 -4.000 991.060 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 1008.230 -4.000 1008.790 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 1025.960 -4.000 1026.520 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met2 ;
        RECT 1043.690 -4.000 1044.250 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 1061.420 -4.000 1061.980 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met2 ;
        RECT 1079.150 -4.000 1079.710 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 1096.880 -4.000 1097.440 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met2 ;
        RECT 1114.610 -4.000 1115.170 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met2 ;
        RECT 1132.340 -4.000 1132.900 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 1150.070 -4.000 1150.630 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 671.360 -4.000 671.920 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met2 ;
        RECT 1167.800 -4.000 1168.360 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 1185.530 -4.000 1186.090 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met2 ;
        RECT 1203.260 -4.000 1203.820 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 1220.990 -4.000 1221.550 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 1238.720 -4.000 1239.280 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 1256.450 -4.000 1257.010 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met2 ;
        RECT 1274.180 -4.000 1274.740 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met2 ;
        RECT 1291.910 -4.000 1292.470 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met2 ;
        RECT 1309.640 -4.000 1310.200 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met2 ;
        RECT 1327.370 -4.000 1327.930 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 689.090 -4.000 689.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 1345.100 -4.000 1345.660 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met2 ;
        RECT 1362.830 -4.000 1363.390 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met2 ;
        RECT 1380.560 -4.000 1381.120 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 1398.290 -4.000 1398.850 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met2 ;
        RECT 1416.020 -4.000 1416.580 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met2 ;
        RECT 1433.750 -4.000 1434.310 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met2 ;
        RECT 1451.480 -4.000 1452.040 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 1469.210 -4.000 1469.770 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met2 ;
        RECT 1486.940 -4.000 1487.500 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 1504.670 -4.000 1505.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 706.820 -4.000 707.380 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met2 ;
        RECT 1522.400 -4.000 1522.960 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met2 ;
        RECT 1540.130 -4.000 1540.690 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met2 ;
        RECT 1557.860 -4.000 1558.420 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 1575.590 -4.000 1576.150 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 1593.320 -4.000 1593.880 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 1611.050 -4.000 1611.610 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 1628.780 -4.000 1629.340 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met2 ;
        RECT 1646.510 -4.000 1647.070 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met2 ;
        RECT 1664.240 -4.000 1664.800 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 1681.970 -4.000 1682.530 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met2 ;
        RECT 724.550 -4.000 725.110 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met2 ;
        RECT 1699.700 -4.000 1700.260 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1717.430 -4.000 1717.990 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1735.160 -4.000 1735.720 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 1752.890 -4.000 1753.450 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 1770.620 -4.000 1771.180 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 1788.350 -4.000 1788.910 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met2 ;
        RECT 1806.080 -4.000 1806.640 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1823.810 -4.000 1824.370 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met2 ;
        RECT 1841.540 -4.000 1842.100 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 1859.270 -4.000 1859.830 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 742.280 -4.000 742.840 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met2 ;
        RECT 1877.000 -4.000 1877.560 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met2 ;
        RECT 1894.730 -4.000 1895.290 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met2 ;
        RECT 1912.460 -4.000 1913.020 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met2 ;
        RECT 1930.190 -4.000 1930.750 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met2 ;
        RECT 1947.920 -4.000 1948.480 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 1965.650 -4.000 1966.210 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met2 ;
        RECT 1983.380 -4.000 1983.940 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met2 ;
        RECT 2001.110 -4.000 2001.670 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 2018.840 -4.000 2019.400 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met2 ;
        RECT 2036.570 -4.000 2037.130 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 760.010 -4.000 760.570 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met2 ;
        RECT 2054.300 -4.000 2054.860 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met2 ;
        RECT 2072.030 -4.000 2072.590 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met2 ;
        RECT 2089.760 -4.000 2090.320 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 2107.490 -4.000 2108.050 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met2 ;
        RECT 2125.220 -4.000 2125.780 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met2 ;
        RECT 2142.950 -4.000 2143.510 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met2 ;
        RECT 2160.680 -4.000 2161.240 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 2178.410 -4.000 2178.970 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met2 ;
        RECT 2196.140 -4.000 2196.700 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 2213.870 -4.000 2214.430 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 777.740 -4.000 778.300 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met2 ;
        RECT 2231.600 -4.000 2232.160 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 2249.330 -4.000 2249.890 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met2 ;
        RECT 2267.060 -4.000 2267.620 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met2 ;
        RECT 2284.790 -4.000 2285.350 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 2302.520 -4.000 2303.080 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met2 ;
        RECT 2320.250 -4.000 2320.810 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 2337.980 -4.000 2338.540 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met2 ;
        RECT 2355.710 -4.000 2356.270 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 2373.440 -4.000 2374.000 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met2 ;
        RECT 2391.170 -4.000 2391.730 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met2 ;
        RECT 795.470 -4.000 796.030 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    PORT
      LAYER met2 ;
        RECT 2893.520 -4.000 2894.080 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    PORT
      LAYER met2 ;
        RECT 2899.430 -4.000 2899.990 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    PORT
      LAYER met2 ;
        RECT 2905.340 -4.000 2905.900 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met2 ;
        RECT 2911.250 -4.000 2911.810 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    PORT
      LAYER met3 ;
        RECT 2911.700 3193.920 2924.000 3217.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2833.630 3143.920 2924.000 3167.920 ;
    END
  END vccd1
  PIN vccd2
    PORT
      LAYER met3 ;
        RECT -14.000 3214.210 -1.700 3238.210 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.000 3164.210 -1.700 3188.210 ;
    END
  END vccd2
  PIN vdda1
    PORT
      LAYER met3 ;
        RECT 2811.595 2697.810 2924.000 2721.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 2747.810 2924.000 2771.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 1171.150 2924.000 1195.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 1121.150 2924.000 1145.150 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met3 ;
        RECT -14.000 1019.440 -1.700 1043.440 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.000 1069.440 -1.700 1093.440 ;
    END
  END vdda2
  PIN vssa1
    PORT
      LAYER met3 ;
        RECT 2597.970 3442.800 2621.970 3514.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2547.970 3442.800 2571.970 3514.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 729.150 2924.000 753.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 679.150 2924.000 703.150 ;
    END
  END vssa1
  PIN vssa2
    PORT
      LAYER met3 ;
        RECT -14.000 2792.210 -1.700 2816.210 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.000 2742.210 -1.700 2766.210 ;
    END
  END vssa2
  PIN vssd1
    PORT
      LAYER met3 ;
        RECT 2883.145 952.150 2924.000 976.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 902.150 2924.000 926.150 ;
    END
  END vssd1
  PIN vssd2
    PORT
      LAYER met3 ;
        RECT -14.000 859.440 -1.700 883.440 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.000 809.440 -1.700 833.440 ;
    END
  END vssd2
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT -2.380 -4.000 -1.820 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 3.530 -4.000 4.090 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 9.440 -4.000 10.000 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 33.080 -4.000 33.640 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 234.020 -4.000 234.580 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 251.750 -4.000 252.310 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 269.480 -4.000 270.040 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 287.210 -4.000 287.770 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 304.940 -4.000 305.500 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 322.670 -4.000 323.230 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 340.400 -4.000 340.960 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 358.130 -4.000 358.690 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 375.860 -4.000 376.420 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 393.590 -4.000 394.150 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 56.720 -4.000 57.280 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 411.320 -4.000 411.880 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 429.050 -4.000 429.610 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 446.780 -4.000 447.340 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 464.510 -4.000 465.070 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 482.240 -4.000 482.800 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 499.970 -4.000 500.530 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 517.700 -4.000 518.260 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 535.430 -4.000 535.990 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 553.160 -4.000 553.720 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 570.890 -4.000 571.450 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 80.360 -4.000 80.920 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 588.620 -4.000 589.180 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 606.350 -4.000 606.910 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 104.000 -4.000 104.560 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 127.640 -4.000 128.200 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 145.370 -4.000 145.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 163.100 -4.000 163.660 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 180.830 -4.000 181.390 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 198.560 -4.000 199.120 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 216.290 -4.000 216.850 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 15.350 -4.000 15.910 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 38.990 -4.000 39.550 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 239.930 -4.000 240.490 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 257.660 -4.000 258.220 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 275.390 -4.000 275.950 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 293.120 -4.000 293.680 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 310.850 -4.000 311.410 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 328.580 -4.000 329.140 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 346.310 -4.000 346.870 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 364.040 -4.000 364.600 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 381.770 -4.000 382.330 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 399.500 -4.000 400.060 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 62.630 -4.000 63.190 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 417.230 -4.000 417.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 434.960 -4.000 435.520 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 452.690 -4.000 453.250 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 470.420 -4.000 470.980 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 488.150 -4.000 488.710 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 505.880 -4.000 506.440 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 523.610 -4.000 524.170 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 541.340 -4.000 541.900 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 559.070 -4.000 559.630 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 576.800 -4.000 577.360 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 86.270 -4.000 86.830 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 594.530 -4.000 595.090 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 612.260 -4.000 612.820 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 109.910 -4.000 110.470 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 133.550 -4.000 134.110 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 151.280 -4.000 151.840 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 169.010 -4.000 169.570 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 186.740 -4.000 187.300 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 204.470 -4.000 205.030 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 222.200 -4.000 222.760 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 44.900 -4.000 45.460 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 245.840 -4.000 246.400 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 263.570 -4.000 264.130 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 281.300 -4.000 281.860 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 299.030 -4.000 299.590 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 316.760 -4.000 317.320 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 334.490 -4.000 335.050 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 352.220 -4.000 352.780 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 369.950 -4.000 370.510 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 387.680 -4.000 388.240 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 405.410 -4.000 405.970 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 68.540 -4.000 69.100 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 423.140 -4.000 423.700 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 440.870 -4.000 441.430 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 458.600 -4.000 459.160 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 476.330 -4.000 476.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 494.060 -4.000 494.620 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 511.790 -4.000 512.350 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 529.520 -4.000 530.080 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 547.250 -4.000 547.810 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 564.980 -4.000 565.540 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 582.710 -4.000 583.270 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 92.180 -4.000 92.740 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 600.440 -4.000 601.000 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 618.170 -4.000 618.730 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 115.820 -4.000 116.380 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 139.460 -4.000 140.020 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 157.190 -4.000 157.750 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 174.920 -4.000 175.480 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 192.650 -4.000 193.210 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 210.380 -4.000 210.940 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 228.110 -4.000 228.670 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 50.810 -4.000 51.370 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 74.450 -4.000 75.010 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 98.090 -4.000 98.650 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 121.730 -4.000 122.290 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 21.260 -4.000 21.820 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 27.170 -4.000 27.730 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 1728.740 3094.200 1855.470 3145.160 ;
      LAYER met1 ;
        RECT 1730.190 3094.210 1853.575 3147.285 ;
      LAYER met2 ;
        RECT 1730.175 3094.205 1853.590 3147.285 ;
      LAYER met3 ;
        RECT 67.030 3452.485 854.070 3471.460 ;
        RECT 865.870 3452.485 866.570 3471.460 ;
        RECT 878.370 3452.650 1112.570 3471.460 ;
        RECT 1124.370 3452.650 1125.070 3471.460 ;
        RECT 1136.870 3452.650 1594.570 3471.460 ;
        RECT 878.370 3452.485 1594.570 3452.650 ;
        RECT 67.030 3247.050 1594.570 3452.485 ;
        RECT 1620.370 3452.565 1621.070 3471.460 ;
        RECT 1632.870 3460.060 1633.570 3471.460 ;
        RECT 1645.370 3460.060 1646.070 3471.460 ;
        RECT 1632.870 3452.565 1646.070 3460.060 ;
        RECT 1620.370 3247.050 1646.070 3452.565 ;
        RECT 1671.870 3452.400 2552.570 3471.460 ;
        RECT 2577.370 3452.400 2602.570 3471.460 ;
        RECT 2627.370 3452.400 2898.095 3471.460 ;
        RECT 1671.870 3422.080 2898.095 3452.400 ;
        RECT 1671.870 3247.050 2552.570 3422.080 ;
        RECT 67.030 3187.405 2552.570 3247.050 ;
        RECT 2577.370 3223.320 2898.095 3422.080 ;
        RECT 2577.370 3198.520 2833.230 3223.320 ;
        RECT 2577.370 3187.405 2898.095 3198.520 ;
        RECT 67.030 3173.320 2898.095 3187.405 ;
        RECT 67.030 3148.520 2833.230 3173.320 ;
        RECT 67.030 2777.210 2898.095 3148.520 ;
        RECT 67.030 2752.410 2811.195 2777.210 ;
        RECT 67.030 2727.210 2898.095 2752.410 ;
        RECT 67.030 2702.410 2811.195 2727.210 ;
        RECT 67.030 2558.610 2898.095 2702.410 ;
        RECT 1700.760 2557.250 2898.095 2558.610 ;
        RECT 67.030 2501.210 2898.095 2557.250 ;
        RECT 67.030 2499.850 2897.695 2501.210 ;
        RECT 67.030 2495.300 2898.095 2499.850 ;
        RECT 67.030 2493.940 2697.070 2495.300 ;
        RECT 67.030 2318.860 2898.095 2493.940 ;
        RECT 1705.795 2317.500 2898.095 2318.860 ;
        RECT 67.030 2312.950 2898.095 2317.500 ;
        RECT 69.885 2311.590 2898.095 2312.950 ;
        RECT 67.030 2279.100 2898.095 2311.590 ;
        RECT 67.030 2277.740 2897.695 2279.100 ;
        RECT 67.030 2273.190 2898.095 2277.740 ;
        RECT 67.030 2271.830 2686.480 2273.190 ;
        RECT 67.030 2102.750 2898.095 2271.830 ;
        RECT 1709.650 2101.390 2898.095 2102.750 ;
        RECT 67.030 2096.840 2898.095 2101.390 ;
        RECT 69.955 2095.480 2898.095 2096.840 ;
        RECT 67.030 2027.440 2898.095 2095.480 ;
        RECT 67.030 2026.080 2667.085 2027.440 ;
        RECT 67.030 981.550 2898.095 2026.080 ;
        RECT 67.030 957.150 86.705 981.550 ;
        RECT 2868.425 957.150 2882.745 981.550 ;
      LAYER met4 ;
        RECT 69.055 955.490 2884.080 3453.685 ;
      LAYER met5 ;
        RECT 1728.910 2985.260 1854.855 3249.955 ;
  END
END DIGITALTBD
END LIBRARY

