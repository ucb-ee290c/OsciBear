VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DIGITALTBD
  CLASS BLOCK ;
  FOREIGN DIGITALTBD ;
  ORIGIN 0.000 0.000 ;
  
  # Reduced from `caravel_user` by (10x10)um (5um per side)
  SIZE 2910.000 BY 3510.000 ;

  PIN VCCD1
    PORT
      LAYER met3 ;
        RECT 2833.630 3198.920 2924.000 3222.920 ;
    END
  END VCCD1
  PIN VDDA1
    PORT
      LAYER met3 ;
        RECT 2811.595 2752.810 2924.000 2776.810 ;
    END
  END VDDA1
  PIN VSSA1
    PORT
      LAYER met3 ;
        RECT 2552.970 3187.805 2576.970 3421.680 ;
    END
  END VSSA1
  PIN VSSD1
    PORT
      LAYER met3 ;
        RECT 87.105 957.150 2868.025 981.150 ;
    END
  END VSSD1
  PIN gpio_analog[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1346.150 2924.000 1346.710 ;
    END
  END gpio_analog[0]
  PIN gpio_analog[10]
    PORT
      LAYER met3 ;
        RECT -4.000 1909.320 2.400 1909.880 ;
    END
  END gpio_analog[10]
  PIN gpio_analog[11]
    PORT
      LAYER met3 ;
        RECT -4.000 1693.210 2.400 1693.770 ;
    END
  END gpio_analog[11]
  PIN gpio_analog[12]
    PORT
      LAYER met3 ;
        RECT -4.000 1477.100 2.400 1477.660 ;
    END
  END gpio_analog[12]
  PIN gpio_analog[13]
    PORT
      LAYER met3 ;
        RECT -4.000 1261.990 2.400 1262.550 ;
    END
  END gpio_analog[13]
  PIN gpio_analog[14]
    PORT
      LAYER met3 ;
        RECT -4.000 623.880 2.400 624.440 ;
    END
  END gpio_analog[14]
  PIN gpio_analog[15]
    PORT
      LAYER met3 ;
        RECT -4.000 407.770 2.400 408.330 ;
    END
  END gpio_analog[15]
  PIN gpio_analog[16]
    PORT
      LAYER met3 ;
        RECT -4.000 191.660 2.400 192.220 ;
    END
  END gpio_analog[16]
  PIN gpio_analog[17]
    PORT
      LAYER met3 ;
        RECT -4.000 84.550 2.400 85.110 ;
    END
  END gpio_analog[17]
  PIN gpio_analog[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1568.260 2924.000 1568.820 ;
    END
  END gpio_analog[1]
  PIN gpio_analog[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1794.370 2924.000 1794.930 ;
    END
  END gpio_analog[2]
  PIN gpio_analog[3]
    PORT
      LAYER met3 ;
        RECT 2667.485 2026.480 2924.000 2027.040 ;
    END
  END gpio_analog[3]
  PIN gpio_analog[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2248.590 2924.000 2249.150 ;
    END
  END gpio_analog[4]
  PIN gpio_analog[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2470.700 2924.000 2471.260 ;
    END
  END gpio_analog[5]
  PIN gpio_analog[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2917.810 2924.000 2918.370 ;
    END
  END gpio_analog[6]
  PIN gpio_analog[7]
    PORT
      LAYER met3 ;
        RECT -4.000 2557.650 1700.360 2558.210 ;
    END
  END gpio_analog[7]
  PIN gpio_analog[8]
    PORT
      LAYER met3 ;
        RECT -4.000 2341.540 2.400 2342.100 ;
    END
  END gpio_analog[8]
  PIN gpio_analog[9]
    PORT
      LAYER met3 ;
        RECT -4.000 2125.430 2.400 2125.990 ;
    END
  END gpio_analog[9]
  PIN gpio_noesd[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 1352.060 2924.000 1352.620 ;
    END
  END gpio_noesd[0]
  PIN gpio_noesd[10]
    PORT
      LAYER met3 ;
        RECT -4.000 1903.410 2.400 1903.970 ;
    END
  END gpio_noesd[10]
  PIN gpio_noesd[11]
    PORT
      LAYER met3 ;
        RECT -4.000 1687.300 2.400 1687.860 ;
    END
  END gpio_noesd[11]
  PIN gpio_noesd[12]
    PORT
      LAYER met3 ;
        RECT -4.000 1471.190 2.400 1471.750 ;
    END
  END gpio_noesd[12]
  PIN gpio_noesd[13]
    PORT
      LAYER met3 ;
        RECT -4.000 1256.080 2.400 1256.640 ;
    END
  END gpio_noesd[13]
  PIN gpio_noesd[14]
    PORT
      LAYER met3 ;
        RECT -4.000 617.970 2.400 618.530 ;
    END
  END gpio_noesd[14]
  PIN gpio_noesd[15]
    PORT
      LAYER met3 ;
        RECT -4.000 401.860 2.400 402.420 ;
    END
  END gpio_noesd[15]
  PIN gpio_noesd[16]
    PORT
      LAYER met3 ;
        RECT -4.000 185.750 2.400 186.310 ;
    END
  END gpio_noesd[16]
  PIN gpio_noesd[17]
    PORT
      LAYER met3 ;
        RECT -4.000 78.640 2.400 79.200 ;
    END
  END gpio_noesd[17]
  PIN gpio_noesd[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 1574.170 2924.000 1574.730 ;
    END
  END gpio_noesd[1]
  PIN gpio_noesd[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1800.280 2924.000 1800.840 ;
    END
  END gpio_noesd[2]
  PIN gpio_noesd[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 2032.390 2924.000 2032.950 ;
    END
  END gpio_noesd[3]
  PIN gpio_noesd[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 2254.500 2924.000 2255.060 ;
    END
  END gpio_noesd[4]
  PIN gpio_noesd[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2476.610 2924.000 2477.170 ;
    END
  END gpio_noesd[5]
  PIN gpio_noesd[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2923.720 2924.000 2924.280 ;
    END
  END gpio_noesd[6]
  PIN gpio_noesd[7]
    PORT
      LAYER met3 ;
        RECT -4.000 2551.740 2.400 2552.300 ;
    END
  END gpio_noesd[7]
  PIN gpio_noesd[8]
    PORT
      LAYER met3 ;
        RECT -4.000 2335.630 2.400 2336.190 ;
    END
  END gpio_noesd[8]
  PIN gpio_noesd[9]
    PORT
      LAYER met3 ;
        RECT -4.000 2119.520 2.400 2120.080 ;
    END
  END gpio_noesd[9]
  PIN io_analog[0]
    PORT
      LAYER met3 ;
        RECT 2911.500 3389.920 2924.000 3414.920 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    PORT
      LAYER met3 ;
        RECT -4.000 3401.210 8.500 3426.210 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    PORT
      LAYER met3 ;
        RECT 2832.970 3511.500 2857.970 3524.000 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    PORT
      LAYER met3 ;
        RECT 2326.970 3511.500 2351.970 3524.000 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    PORT
      LAYER met3 ;
        RECT 2066.970 3511.500 2091.970 3524.000 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    PORT
      LAYER met3 ;
        RECT 1646.470 3247.450 1671.470 3524.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1594.970 3247.450 1619.970 3524.000 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    PORT
      LAYER met3 ;
        RECT 1137.970 3511.500 1162.970 3524.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1086.470 3511.500 1111.470 3524.000 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    PORT
      LAYER met3 ;
        RECT 879.470 3511.500 904.470 3524.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 827.970 3511.500 852.970 3524.000 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    PORT
      LAYER met3 ;
        RECT 600.970 3511.500 625.970 3524.000 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    PORT
      LAYER met3 ;
        RECT 340.970 3511.500 365.970 3524.000 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    PORT
      LAYER met3 ;
        RECT 80.970 3511.500 105.970 3524.000 ;
    END
  END io_analog[9]
  PIN io_clamp_high[0]
    PORT
      LAYER met3 ;
        RECT 1633.970 3460.460 1644.970 3524.000 ;
    END
  END io_clamp_high[0]
  PIN io_clamp_high[1]
    PORT
      LAYER met3 ;
        RECT 1125.470 3453.050 1136.470 3524.000 ;
    END
  END io_clamp_high[1]
  PIN io_clamp_high[2]
    PORT
      LAYER met3 ;
        RECT 866.970 3452.885 877.970 3524.000 ;
    END
  END io_clamp_high[2]
  PIN io_clamp_low[0]
    PORT
      LAYER met3 ;
        RECT 1621.470 3452.965 1632.470 3524.000 ;
    END
  END io_clamp_low[0]
  PIN io_clamp_low[1]
    PORT
      LAYER met3 ;
        RECT 1112.970 3453.050 1123.970 3524.000 ;
    END
  END io_clamp_low[1]
  PIN io_clamp_low[2]
    PORT
      LAYER met3 ;
        RECT 854.470 3452.885 865.470 3524.000 ;
    END
  END io_clamp_low[2]
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 13.630 2924.000 14.190 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2044.210 2924.000 2044.770 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2266.320 2924.000 2266.880 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2488.430 2924.000 2488.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2935.540 2924.000 2936.100 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met3 ;
        RECT -4.000 2539.920 2.400 2540.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met3 ;
        RECT -4.000 2323.810 2.400 2324.370 ;
    END
  END io_in[15]
  PIN io_in[16]
    PORT
      LAYER met3 ;
        RECT -4.000 2107.700 2.400 2108.260 ;
    END
  END io_in[16]
  PIN io_in[17]
    PORT
      LAYER met3 ;
        RECT -4.000 1891.590 2.400 1892.150 ;
    END
  END io_in[17]
  PIN io_in[18]
    PORT
      LAYER met3 ;
        RECT -4.000 1675.480 2.400 1676.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    PORT
      LAYER met3 ;
        RECT -4.000 1459.370 2.400 1459.930 ;
    END
  END io_in[19]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 37.270 2924.000 37.830 ;
    END
  END io_in[1]
  PIN io_in[20]
    PORT
      LAYER met3 ;
        RECT -4.000 1244.260 2.400 1244.820 ;
    END
  END io_in[20]
  PIN io_in[21]
    PORT
      LAYER met3 ;
        RECT -4.000 606.150 2.400 606.710 ;
    END
  END io_in[21]
  PIN io_in[22]
    PORT
      LAYER met3 ;
        RECT -4.000 390.040 2.400 390.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    PORT
      LAYER met3 ;
        RECT -4.000 173.930 2.400 174.490 ;
    END
  END io_in[23]
  PIN io_in[24]
    PORT
      LAYER met3 ;
        RECT -4.000 66.820 2.400 67.380 ;
    END
  END io_in[24]
  PIN io_in[25]
    PORT
      LAYER met3 ;
        RECT -4.000 43.180 2.400 43.740 ;
    END
  END io_in[25]
  PIN io_in[26]
    PORT
      LAYER met3 ;
        RECT -4.000 19.540 2.400 20.100 ;
    END
  END io_in[26]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 60.910 2924.000 61.470 ;
    END
  END io_in[2]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 84.550 2924.000 85.110 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 108.190 2924.000 108.750 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 240.480 2924.000 241.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 463.770 2924.000 464.330 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1363.880 2924.000 1364.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1585.990 2924.000 1586.550 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1812.100 2924.000 1812.660 ;
    END
  END io_in[9]
  PIN io_in_3v3[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 7.720 2924.000 8.280 ;
    END
  END io_in_3v3[0]
  PIN io_in_3v3[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2038.300 2924.000 2038.860 ;
    END
  END io_in_3v3[10]
  PIN io_in_3v3[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 2260.410 2924.000 2260.970 ;
    END
  END io_in_3v3[11]
  PIN io_in_3v3[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 2482.520 2924.000 2483.080 ;
    END
  END io_in_3v3[12]
  PIN io_in_3v3[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2929.630 2924.000 2930.190 ;
    END
  END io_in_3v3[13]
  PIN io_in_3v3[14]
    PORT
      LAYER met3 ;
        RECT -4.000 2545.830 2.400 2546.390 ;
    END
  END io_in_3v3[14]
  PIN io_in_3v3[15]
    PORT
      LAYER met3 ;
        RECT -4.000 2329.720 2.400 2330.280 ;
    END
  END io_in_3v3[15]
  PIN io_in_3v3[16]
    PORT
      LAYER met3 ;
        RECT -4.000 2113.610 2.400 2114.170 ;
    END
  END io_in_3v3[16]
  PIN io_in_3v3[17]
    PORT
      LAYER met3 ;
        RECT -4.000 1897.500 2.400 1898.060 ;
    END
  END io_in_3v3[17]
  PIN io_in_3v3[18]
    PORT
      LAYER met3 ;
        RECT -4.000 1681.390 2.400 1681.950 ;
    END
  END io_in_3v3[18]
  PIN io_in_3v3[19]
    PORT
      LAYER met3 ;
        RECT -4.000 1465.280 2.400 1465.840 ;
    END
  END io_in_3v3[19]
  PIN io_in_3v3[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 31.360 2924.000 31.920 ;
    END
  END io_in_3v3[1]
  PIN io_in_3v3[20]
    PORT
      LAYER met3 ;
        RECT -4.000 1250.170 2.400 1250.730 ;
    END
  END io_in_3v3[20]
  PIN io_in_3v3[21]
    PORT
      LAYER met3 ;
        RECT -4.000 612.060 2.400 612.620 ;
    END
  END io_in_3v3[21]
  PIN io_in_3v3[22]
    PORT
      LAYER met3 ;
        RECT -4.000 395.950 2.400 396.510 ;
    END
  END io_in_3v3[22]
  PIN io_in_3v3[23]
    PORT
      LAYER met3 ;
        RECT -4.000 179.840 2.400 180.400 ;
    END
  END io_in_3v3[23]
  PIN io_in_3v3[24]
    PORT
      LAYER met3 ;
        RECT -4.000 72.730 2.400 73.290 ;
    END
  END io_in_3v3[24]
  PIN io_in_3v3[25]
    PORT
      LAYER met3 ;
        RECT -4.000 49.090 2.400 49.650 ;
    END
  END io_in_3v3[25]
  PIN io_in_3v3[26]
    PORT
      LAYER met3 ;
        RECT -4.000 25.450 2.400 26.010 ;
    END
  END io_in_3v3[26]
  PIN io_in_3v3[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 55.000 2924.000 55.560 ;
    END
  END io_in_3v3[2]
  PIN io_in_3v3[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 78.640 2924.000 79.200 ;
    END
  END io_in_3v3[3]
  PIN io_in_3v3[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 102.280 2924.000 102.840 ;
    END
  END io_in_3v3[4]
  PIN io_in_3v3[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 234.570 2924.000 235.130 ;
    END
  END io_in_3v3[5]
  PIN io_in_3v3[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 457.860 2924.000 458.420 ;
    END
  END io_in_3v3[6]
  PIN io_in_3v3[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1357.970 2924.000 1358.530 ;
    END
  END io_in_3v3[7]
  PIN io_in_3v3[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1580.080 2924.000 1580.640 ;
    END
  END io_in_3v3[8]
  PIN io_in_3v3[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1806.190 2924.000 1806.750 ;
    END
  END io_in_3v3[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 25.450 2924.000 26.010 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2056.030 2924.000 2056.590 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met3 ;
        RECT 2898.095 2278.140 2924.000 2278.700 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met3 ;
        RECT 2898.095 2500.250 2924.000 2500.810 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2947.360 2924.000 2947.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT -4.000 2528.100 2.400 2528.660 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met3 ;
        RECT -4.000 2311.990 69.485 2312.550 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    PORT
      LAYER met3 ;
        RECT -4.000 2095.880 69.555 2096.440 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    PORT
      LAYER met3 ;
        RECT -4.000 1879.770 2.400 1880.330 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    PORT
      LAYER met3 ;
        RECT -4.000 1663.660 2.400 1664.220 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    PORT
      LAYER met3 ;
        RECT -4.000 1447.550 2.400 1448.110 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 49.090 2924.000 49.650 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    PORT
      LAYER met3 ;
        RECT -4.000 1232.440 2.400 1233.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    PORT
      LAYER met3 ;
        RECT -4.000 594.330 2.400 594.890 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    PORT
      LAYER met3 ;
        RECT -4.000 378.220 2.400 378.780 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    PORT
      LAYER met3 ;
        RECT -4.000 162.110 2.400 162.670 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    PORT
      LAYER met3 ;
        RECT -4.000 55.000 2.400 55.560 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    PORT
      LAYER met3 ;
        RECT -4.000 31.360 2.400 31.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    PORT
      LAYER met3 ;
        RECT -4.000 7.720 2.400 8.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 72.730 2924.000 73.290 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 96.370 2924.000 96.930 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 120.010 2924.000 120.570 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 252.300 2924.000 252.860 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 475.590 2924.000 476.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1375.700 2924.000 1376.260 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1597.810 2924.000 1598.370 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1823.920 2924.000 1824.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 19.540 2924.000 20.100 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2050.120 2924.000 2050.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 2686.880 2272.230 2924.000 2272.790 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT 2697.470 2494.340 2924.000 2494.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2941.450 2924.000 2942.010 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met3 ;
        RECT -4.000 2534.010 2.400 2534.570 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met3 ;
        RECT -4.000 2317.900 1705.395 2318.460 ;
    END
  END io_out[15]
  PIN io_out[16]
    PORT
      LAYER met3 ;
        RECT -4.000 2101.790 1709.250 2102.350 ;
    END
  END io_out[16]
  PIN io_out[17]
    PORT
      LAYER met3 ;
        RECT -4.000 1885.680 2.400 1886.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    PORT
      LAYER met3 ;
        RECT -4.000 1669.570 2.400 1670.130 ;
    END
  END io_out[18]
  PIN io_out[19]
    PORT
      LAYER met3 ;
        RECT -4.000 1453.460 2.400 1454.020 ;
    END
  END io_out[19]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 43.180 2924.000 43.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    PORT
      LAYER met3 ;
        RECT -4.000 1238.350 2.400 1238.910 ;
    END
  END io_out[20]
  PIN io_out[21]
    PORT
      LAYER met3 ;
        RECT -4.000 600.240 2.400 600.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    PORT
      LAYER met3 ;
        RECT -4.000 384.130 2.400 384.690 ;
    END
  END io_out[22]
  PIN io_out[23]
    PORT
      LAYER met3 ;
        RECT -4.000 168.020 2.400 168.580 ;
    END
  END io_out[23]
  PIN io_out[24]
    PORT
      LAYER met3 ;
        RECT -4.000 60.910 2.400 61.470 ;
    END
  END io_out[24]
  PIN io_out[25]
    PORT
      LAYER met3 ;
        RECT -4.000 37.270 2.400 37.830 ;
    END
  END io_out[25]
  PIN io_out[26]
    PORT
      LAYER met3 ;
        RECT -4.000 13.630 2.400 14.190 ;
    END
  END io_out[26]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 66.820 2924.000 67.380 ;
    END
  END io_out[2]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 90.460 2924.000 91.020 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 114.100 2924.000 114.660 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 246.390 2924.000 246.950 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 469.680 2924.000 470.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 1369.790 2924.000 1370.350 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 1591.900 2924.000 1592.460 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1818.010 2924.000 1818.570 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 629.080 -4.000 629.640 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met2 ;
        RECT 2402.080 -4.000 2402.640 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met2 ;
        RECT 2419.810 -4.000 2420.370 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 2437.540 -4.000 2438.100 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met2 ;
        RECT 2455.270 -4.000 2455.830 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met2 ;
        RECT 2473.000 -4.000 2473.560 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 2490.730 -4.000 2491.290 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 2508.460 -4.000 2509.020 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met2 ;
        RECT 2526.190 -4.000 2526.750 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met2 ;
        RECT 2543.920 -4.000 2544.480 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met2 ;
        RECT 2561.650 -4.000 2562.210 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met2 ;
        RECT 806.380 -4.000 806.940 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met2 ;
        RECT 2579.380 -4.000 2579.940 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met2 ;
        RECT 2597.110 -4.000 2597.670 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met2 ;
        RECT 2614.840 -4.000 2615.400 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met2 ;
        RECT 2632.570 -4.000 2633.130 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met2 ;
        RECT 2650.300 -4.000 2650.860 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 2668.030 -4.000 2668.590 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 2685.760 -4.000 2686.320 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met2 ;
        RECT 2703.490 -4.000 2704.050 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met2 ;
        RECT 2721.220 -4.000 2721.780 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met2 ;
        RECT 2738.950 -4.000 2739.510 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 824.110 -4.000 824.670 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met2 ;
        RECT 2756.680 -4.000 2757.240 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 2774.410 -4.000 2774.970 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 2792.140 -4.000 2792.700 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met2 ;
        RECT 2809.870 -4.000 2810.430 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 2827.600 -4.000 2828.160 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 2845.330 -4.000 2845.890 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met2 ;
        RECT 2863.060 -4.000 2863.620 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2880.790 -4.000 2881.350 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met2 ;
        RECT 841.840 -4.000 842.400 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met2 ;
        RECT 859.570 -4.000 860.130 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met2 ;
        RECT 877.300 -4.000 877.860 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met2 ;
        RECT 895.030 -4.000 895.590 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met2 ;
        RECT 912.760 -4.000 913.320 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met2 ;
        RECT 930.490 -4.000 931.050 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met2 ;
        RECT 948.220 -4.000 948.780 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 965.950 -4.000 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 646.810 -4.000 647.370 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met2 ;
        RECT 983.680 -4.000 984.240 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 1001.410 -4.000 1001.970 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 1019.140 -4.000 1019.700 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met2 ;
        RECT 1036.870 -4.000 1037.430 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met2 ;
        RECT 1054.600 -4.000 1055.160 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 1072.330 -4.000 1072.890 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 1090.060 -4.000 1090.620 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 1107.790 -4.000 1108.350 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met2 ;
        RECT 1125.520 -4.000 1126.080 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met2 ;
        RECT 1143.250 -4.000 1143.810 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 664.540 -4.000 665.100 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met2 ;
        RECT 1160.980 -4.000 1161.540 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met2 ;
        RECT 1178.710 -4.000 1179.270 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 1196.440 -4.000 1197.000 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met2 ;
        RECT 1214.170 -4.000 1214.730 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met2 ;
        RECT 1231.900 -4.000 1232.460 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met2 ;
        RECT 1249.630 -4.000 1250.190 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 1267.360 -4.000 1267.920 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 1285.090 -4.000 1285.650 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 1302.820 -4.000 1303.380 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 1320.550 -4.000 1321.110 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met2 ;
        RECT 682.270 -4.000 682.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 1338.280 -4.000 1338.840 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met2 ;
        RECT 1356.010 -4.000 1356.570 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met2 ;
        RECT 1373.740 -4.000 1374.300 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met2 ;
        RECT 1391.470 -4.000 1392.030 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met2 ;
        RECT 1409.200 -4.000 1409.760 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 1426.930 -4.000 1427.490 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 1444.660 -4.000 1445.220 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met2 ;
        RECT 1462.390 -4.000 1462.950 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met2 ;
        RECT 1480.120 -4.000 1480.680 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met2 ;
        RECT 1497.850 -4.000 1498.410 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 700.000 -4.000 700.560 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 1515.580 -4.000 1516.140 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met2 ;
        RECT 1533.310 -4.000 1533.870 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met2 ;
        RECT 1551.040 -4.000 1551.600 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 1568.770 -4.000 1569.330 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 1586.500 -4.000 1587.060 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met2 ;
        RECT 1604.230 -4.000 1604.790 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met2 ;
        RECT 1621.960 -4.000 1622.520 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met2 ;
        RECT 1639.690 -4.000 1640.250 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 1657.420 -4.000 1657.980 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met2 ;
        RECT 1675.150 -4.000 1675.710 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met2 ;
        RECT 717.730 -4.000 718.290 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 1692.880 -4.000 1693.440 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 1710.610 -4.000 1711.170 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met2 ;
        RECT 1728.340 -4.000 1728.900 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met2 ;
        RECT 1746.070 -4.000 1746.630 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met2 ;
        RECT 1763.800 -4.000 1764.360 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.000 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met2 ;
        RECT 1799.260 -4.000 1799.820 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 1816.990 -4.000 1817.550 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met2 ;
        RECT 1834.720 -4.000 1835.280 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met2 ;
        RECT 1852.450 -4.000 1853.010 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met2 ;
        RECT 735.460 -4.000 736.020 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met2 ;
        RECT 1870.180 -4.000 1870.740 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met2 ;
        RECT 1887.910 -4.000 1888.470 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 1905.640 -4.000 1906.200 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met2 ;
        RECT 1923.370 -4.000 1923.930 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met2 ;
        RECT 1941.100 -4.000 1941.660 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 1958.830 -4.000 1959.390 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met2 ;
        RECT 1976.560 -4.000 1977.120 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 1994.290 -4.000 1994.850 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 2012.020 -4.000 2012.580 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met2 ;
        RECT 2029.750 -4.000 2030.310 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 753.190 -4.000 753.750 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met2 ;
        RECT 2047.480 -4.000 2048.040 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 2065.210 -4.000 2065.770 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 2082.940 -4.000 2083.500 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met2 ;
        RECT 2100.670 -4.000 2101.230 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met2 ;
        RECT 2118.400 -4.000 2118.960 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met2 ;
        RECT 2136.130 -4.000 2136.690 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met2 ;
        RECT 2153.860 -4.000 2154.420 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 2171.590 -4.000 2172.150 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met2 ;
        RECT 2189.320 -4.000 2189.880 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 2207.050 -4.000 2207.610 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 770.920 -4.000 771.480 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met2 ;
        RECT 2224.780 -4.000 2225.340 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met2 ;
        RECT 2242.510 -4.000 2243.070 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met2 ;
        RECT 2260.240 -4.000 2260.800 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met2 ;
        RECT 2277.970 -4.000 2278.530 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met2 ;
        RECT 2295.700 -4.000 2296.260 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met2 ;
        RECT 2313.430 -4.000 2313.990 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met2 ;
        RECT 2331.160 -4.000 2331.720 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met2 ;
        RECT 2348.890 -4.000 2349.450 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 2366.620 -4.000 2367.180 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met2 ;
        RECT 2384.350 -4.000 2384.910 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 788.650 -4.000 789.210 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met2 ;
        RECT 634.990 -4.000 635.550 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 2407.990 -4.000 2408.550 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 2425.720 -4.000 2426.280 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 2443.450 -4.000 2444.010 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met2 ;
        RECT 2461.180 -4.000 2461.740 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 2478.910 -4.000 2479.470 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met2 ;
        RECT 2496.640 -4.000 2497.200 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 2514.370 -4.000 2514.930 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met2 ;
        RECT 2532.100 -4.000 2532.660 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met2 ;
        RECT 2549.830 -4.000 2550.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 2567.560 -4.000 2568.120 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met2 ;
        RECT 812.290 -4.000 812.850 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met2 ;
        RECT 2585.290 -4.000 2585.850 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met2 ;
        RECT 2603.020 -4.000 2603.580 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met2 ;
        RECT 2620.750 -4.000 2621.310 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 2638.480 -4.000 2639.040 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 2656.210 -4.000 2656.770 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 2673.940 -4.000 2674.500 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 2691.670 -4.000 2692.230 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met2 ;
        RECT 2709.400 -4.000 2709.960 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met2 ;
        RECT 2727.130 -4.000 2727.690 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met2 ;
        RECT 2744.860 -4.000 2745.420 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 830.020 -4.000 830.580 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 2762.590 -4.000 2763.150 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 2780.320 -4.000 2780.880 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 2798.050 -4.000 2798.610 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met2 ;
        RECT 2815.780 -4.000 2816.340 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met2 ;
        RECT 2833.510 -4.000 2834.070 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met2 ;
        RECT 2851.240 -4.000 2851.800 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.000 2869.530 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met2 ;
        RECT 2886.700 -4.000 2887.260 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 847.750 -4.000 848.310 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met2 ;
        RECT 865.480 -4.000 866.040 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met2 ;
        RECT 883.210 -4.000 883.770 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met2 ;
        RECT 900.940 -4.000 901.500 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 918.670 -4.000 919.230 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met2 ;
        RECT 936.400 -4.000 936.960 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 954.130 -4.000 954.690 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 971.860 -4.000 972.420 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met2 ;
        RECT 652.720 -4.000 653.280 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met2 ;
        RECT 989.590 -4.000 990.150 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met2 ;
        RECT 1007.320 -4.000 1007.880 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met2 ;
        RECT 1025.050 -4.000 1025.610 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met2 ;
        RECT 1042.780 -4.000 1043.340 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met2 ;
        RECT 1060.510 -4.000 1061.070 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 1078.240 -4.000 1078.800 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met2 ;
        RECT 1095.970 -4.000 1096.530 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met2 ;
        RECT 1113.700 -4.000 1114.260 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 1131.430 -4.000 1131.990 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 1149.160 -4.000 1149.720 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 670.450 -4.000 671.010 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 1166.890 -4.000 1167.450 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met2 ;
        RECT 1184.620 -4.000 1185.180 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met2 ;
        RECT 1202.350 -4.000 1202.910 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met2 ;
        RECT 1220.080 -4.000 1220.640 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.000 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met2 ;
        RECT 1255.540 -4.000 1256.100 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 1273.270 -4.000 1273.830 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met2 ;
        RECT 1291.000 -4.000 1291.560 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met2 ;
        RECT 1308.730 -4.000 1309.290 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met2 ;
        RECT 1326.460 -4.000 1327.020 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met2 ;
        RECT 688.180 -4.000 688.740 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met2 ;
        RECT 1344.190 -4.000 1344.750 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 1361.920 -4.000 1362.480 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 1379.650 -4.000 1380.210 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met2 ;
        RECT 1397.380 -4.000 1397.940 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 1415.110 -4.000 1415.670 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 1432.840 -4.000 1433.400 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 1450.570 -4.000 1451.130 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met2 ;
        RECT 1468.300 -4.000 1468.860 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 1486.030 -4.000 1486.590 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 1503.760 -4.000 1504.320 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 705.910 -4.000 706.470 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met2 ;
        RECT 1521.490 -4.000 1522.050 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 1539.220 -4.000 1539.780 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met2 ;
        RECT 1556.950 -4.000 1557.510 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 1574.680 -4.000 1575.240 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 1592.410 -4.000 1592.970 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met2 ;
        RECT 1610.140 -4.000 1610.700 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 1627.870 -4.000 1628.430 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 1645.600 -4.000 1646.160 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met2 ;
        RECT 1663.330 -4.000 1663.890 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met2 ;
        RECT 1681.060 -4.000 1681.620 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 723.640 -4.000 724.200 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met2 ;
        RECT 1698.790 -4.000 1699.350 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met2 ;
        RECT 1716.520 -4.000 1717.080 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1734.250 -4.000 1734.810 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 1751.980 -4.000 1752.540 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met2 ;
        RECT 1769.710 -4.000 1770.270 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 1787.440 -4.000 1788.000 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met2 ;
        RECT 1805.170 -4.000 1805.730 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met2 ;
        RECT 1822.900 -4.000 1823.460 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met2 ;
        RECT 1840.630 -4.000 1841.190 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met2 ;
        RECT 1858.360 -4.000 1858.920 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 741.370 -4.000 741.930 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 1876.090 -4.000 1876.650 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met2 ;
        RECT 1893.820 -4.000 1894.380 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 1911.550 -4.000 1912.110 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1929.280 -4.000 1929.840 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 1947.010 -4.000 1947.570 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 1964.740 -4.000 1965.300 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met2 ;
        RECT 1982.470 -4.000 1983.030 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met2 ;
        RECT 2000.200 -4.000 2000.760 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 2017.930 -4.000 2018.490 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met2 ;
        RECT 2035.660 -4.000 2036.220 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met2 ;
        RECT 759.100 -4.000 759.660 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met2 ;
        RECT 2053.390 -4.000 2053.950 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met2 ;
        RECT 2071.120 -4.000 2071.680 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 2088.850 -4.000 2089.410 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met2 ;
        RECT 2106.580 -4.000 2107.140 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 2124.310 -4.000 2124.870 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 2142.040 -4.000 2142.600 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 2159.770 -4.000 2160.330 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 2177.500 -4.000 2178.060 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met2 ;
        RECT 2195.230 -4.000 2195.790 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met2 ;
        RECT 2212.960 -4.000 2213.520 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met2 ;
        RECT 776.830 -4.000 777.390 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 2230.690 -4.000 2231.250 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 2248.420 -4.000 2248.980 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 2266.150 -4.000 2266.710 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 2283.880 -4.000 2284.440 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 2301.610 -4.000 2302.170 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met2 ;
        RECT 2319.340 -4.000 2319.900 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 2337.070 -4.000 2337.630 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 2354.800 -4.000 2355.360 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 2372.530 -4.000 2373.090 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 2390.260 -4.000 2390.820 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met2 ;
        RECT 794.560 -4.000 795.120 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 640.900 -4.000 641.460 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met2 ;
        RECT 2413.900 -4.000 2414.460 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met2 ;
        RECT 2431.630 -4.000 2432.190 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 2449.360 -4.000 2449.920 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 2467.090 -4.000 2467.650 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 2484.820 -4.000 2485.380 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met2 ;
        RECT 2502.550 -4.000 2503.110 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 2520.280 -4.000 2520.840 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 2538.010 -4.000 2538.570 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met2 ;
        RECT 2555.740 -4.000 2556.300 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 2573.470 -4.000 2574.030 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 818.200 -4.000 818.760 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 2591.200 -4.000 2591.760 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 2608.930 -4.000 2609.490 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met2 ;
        RECT 2626.660 -4.000 2627.220 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 2644.390 -4.000 2644.950 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met2 ;
        RECT 2662.120 -4.000 2662.680 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 2679.850 -4.000 2680.410 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met2 ;
        RECT 2697.580 -4.000 2698.140 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 2715.310 -4.000 2715.870 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 2733.040 -4.000 2733.600 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met2 ;
        RECT 2750.770 -4.000 2751.330 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 835.930 -4.000 836.490 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 2768.500 -4.000 2769.060 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met2 ;
        RECT 2786.230 -4.000 2786.790 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met2 ;
        RECT 2803.960 -4.000 2804.520 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 2821.690 -4.000 2822.250 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 2839.420 -4.000 2839.980 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 2857.150 -4.000 2857.710 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 2874.880 -4.000 2875.440 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met2 ;
        RECT 2892.610 -4.000 2893.170 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met2 ;
        RECT 853.660 -4.000 854.220 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met2 ;
        RECT 871.390 -4.000 871.950 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met2 ;
        RECT 889.120 -4.000 889.680 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met2 ;
        RECT 906.850 -4.000 907.410 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met2 ;
        RECT 924.580 -4.000 925.140 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 942.310 -4.000 942.870 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met2 ;
        RECT 960.040 -4.000 960.600 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met2 ;
        RECT 977.770 -4.000 978.330 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 658.630 -4.000 659.190 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met2 ;
        RECT 995.500 -4.000 996.060 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 1013.230 -4.000 1013.790 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 1030.960 -4.000 1031.520 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met2 ;
        RECT 1048.690 -4.000 1049.250 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 1066.420 -4.000 1066.980 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met2 ;
        RECT 1084.150 -4.000 1084.710 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 1101.880 -4.000 1102.440 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met2 ;
        RECT 1119.610 -4.000 1120.170 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met2 ;
        RECT 1137.340 -4.000 1137.900 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 1155.070 -4.000 1155.630 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 676.360 -4.000 676.920 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met2 ;
        RECT 1172.800 -4.000 1173.360 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 1190.530 -4.000 1191.090 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met2 ;
        RECT 1208.260 -4.000 1208.820 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 1225.990 -4.000 1226.550 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 1243.720 -4.000 1244.280 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 1261.450 -4.000 1262.010 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met2 ;
        RECT 1279.180 -4.000 1279.740 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met2 ;
        RECT 1296.910 -4.000 1297.470 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met2 ;
        RECT 1314.640 -4.000 1315.200 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met2 ;
        RECT 1332.370 -4.000 1332.930 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 694.090 -4.000 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 1350.100 -4.000 1350.660 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met2 ;
        RECT 1367.830 -4.000 1368.390 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met2 ;
        RECT 1385.560 -4.000 1386.120 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 1403.290 -4.000 1403.850 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met2 ;
        RECT 1421.020 -4.000 1421.580 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met2 ;
        RECT 1438.750 -4.000 1439.310 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met2 ;
        RECT 1456.480 -4.000 1457.040 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 1474.210 -4.000 1474.770 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met2 ;
        RECT 1491.940 -4.000 1492.500 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.000 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 711.820 -4.000 712.380 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met2 ;
        RECT 1527.400 -4.000 1527.960 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met2 ;
        RECT 1545.130 -4.000 1545.690 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met2 ;
        RECT 1562.860 -4.000 1563.420 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 1580.590 -4.000 1581.150 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 1598.320 -4.000 1598.880 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 1616.050 -4.000 1616.610 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 1633.780 -4.000 1634.340 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met2 ;
        RECT 1651.510 -4.000 1652.070 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met2 ;
        RECT 1669.240 -4.000 1669.800 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 1686.970 -4.000 1687.530 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met2 ;
        RECT 729.550 -4.000 730.110 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met2 ;
        RECT 1704.700 -4.000 1705.260 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1722.430 -4.000 1722.990 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1740.160 -4.000 1740.720 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 1757.890 -4.000 1758.450 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 1775.620 -4.000 1776.180 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 1793.350 -4.000 1793.910 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met2 ;
        RECT 1811.080 -4.000 1811.640 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1828.810 -4.000 1829.370 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met2 ;
        RECT 1846.540 -4.000 1847.100 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 1864.270 -4.000 1864.830 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 747.280 -4.000 747.840 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met2 ;
        RECT 1882.000 -4.000 1882.560 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met2 ;
        RECT 1899.730 -4.000 1900.290 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met2 ;
        RECT 1917.460 -4.000 1918.020 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met2 ;
        RECT 1935.190 -4.000 1935.750 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met2 ;
        RECT 1952.920 -4.000 1953.480 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 1970.650 -4.000 1971.210 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met2 ;
        RECT 1988.380 -4.000 1988.940 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met2 ;
        RECT 2006.110 -4.000 2006.670 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 2023.840 -4.000 2024.400 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met2 ;
        RECT 2041.570 -4.000 2042.130 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 765.010 -4.000 765.570 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met2 ;
        RECT 2059.300 -4.000 2059.860 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met2 ;
        RECT 2077.030 -4.000 2077.590 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met2 ;
        RECT 2094.760 -4.000 2095.320 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 2112.490 -4.000 2113.050 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met2 ;
        RECT 2130.220 -4.000 2130.780 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met2 ;
        RECT 2147.950 -4.000 2148.510 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met2 ;
        RECT 2165.680 -4.000 2166.240 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 2183.410 -4.000 2183.970 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met2 ;
        RECT 2201.140 -4.000 2201.700 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 2218.870 -4.000 2219.430 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 782.740 -4.000 783.300 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met2 ;
        RECT 2236.600 -4.000 2237.160 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 2254.330 -4.000 2254.890 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met2 ;
        RECT 2272.060 -4.000 2272.620 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met2 ;
        RECT 2289.790 -4.000 2290.350 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 2307.520 -4.000 2308.080 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met2 ;
        RECT 2325.250 -4.000 2325.810 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 2342.980 -4.000 2343.540 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met2 ;
        RECT 2360.710 -4.000 2361.270 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 2378.440 -4.000 2379.000 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met2 ;
        RECT 2396.170 -4.000 2396.730 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met2 ;
        RECT 800.470 -4.000 801.030 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    PORT
      LAYER met2 ;
        RECT 2898.520 -4.000 2899.080 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    PORT
      LAYER met2 ;
        RECT 2904.430 -4.000 2904.990 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    PORT
      LAYER met2 ;
        RECT 2910.340 -4.000 2910.900 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met2 ;
        RECT 2916.250 -4.000 2916.810 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    PORT
      LAYER met3 ;
        RECT 2911.700 3198.920 2924.000 3222.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2833.630 3148.920 2924.000 3172.920 ;
    END
  END vccd1
  PIN vccd2
    PORT
      LAYER met3 ;
        RECT -4.000 3219.210 8.300 3243.210 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.000 3169.210 8.300 3193.210 ;
    END
  END vccd2
  PIN vdda1
    PORT
      LAYER met3 ;
        RECT 2811.595 2702.810 2924.000 2726.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 2752.810 2924.000 2776.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 1176.150 2924.000 1200.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 1126.150 2924.000 1150.150 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met3 ;
        RECT -4.000 1024.440 8.300 1048.440 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.000 1074.440 8.300 1098.440 ;
    END
  END vdda2
  PIN vssa1
    PORT
      LAYER met3 ;
        RECT 2602.970 3452.800 2626.970 3524.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2552.970 3452.800 2576.970 3524.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 734.150 2924.000 758.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 684.150 2924.000 708.150 ;
    END
  END vssa1
  PIN vssa2
    PORT
      LAYER met3 ;
        RECT -4.000 2797.210 8.300 2821.210 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.000 2747.210 8.300 2771.210 ;
    END
  END vssa2
  PIN vssd1
    PORT
      LAYER met3 ;
        RECT 2883.145 957.150 2924.000 981.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 2911.700 907.150 2924.000 931.150 ;
    END
  END vssd1
  PIN vssd2
    PORT
      LAYER met3 ;
        RECT -4.000 864.440 8.300 888.440 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.000 814.440 8.300 838.440 ;
    END
  END vssd2
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 2.620 -4.000 3.180 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 8.530 -4.000 9.090 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 14.440 -4.000 15.000 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 38.080 -4.000 38.640 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 239.020 -4.000 239.580 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 256.750 -4.000 257.310 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 274.480 -4.000 275.040 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 292.210 -4.000 292.770 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 309.940 -4.000 310.500 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 327.670 -4.000 328.230 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 345.400 -4.000 345.960 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 363.130 -4.000 363.690 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 380.860 -4.000 381.420 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 398.590 -4.000 399.150 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 61.720 -4.000 62.280 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 416.320 -4.000 416.880 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 434.050 -4.000 434.610 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 451.780 -4.000 452.340 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 469.510 -4.000 470.070 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 487.240 -4.000 487.800 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 504.970 -4.000 505.530 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 522.700 -4.000 523.260 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 540.430 -4.000 540.990 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 558.160 -4.000 558.720 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 575.890 -4.000 576.450 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 85.360 -4.000 85.920 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 593.620 -4.000 594.180 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 611.350 -4.000 611.910 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 109.000 -4.000 109.560 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 132.640 -4.000 133.200 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 150.370 -4.000 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 168.100 -4.000 168.660 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 185.830 -4.000 186.390 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 203.560 -4.000 204.120 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 221.290 -4.000 221.850 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 20.350 -4.000 20.910 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 43.990 -4.000 44.550 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 244.930 -4.000 245.490 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 262.660 -4.000 263.220 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 280.390 -4.000 280.950 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 298.120 -4.000 298.680 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 315.850 -4.000 316.410 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 333.580 -4.000 334.140 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 351.310 -4.000 351.870 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 369.040 -4.000 369.600 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 386.770 -4.000 387.330 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 404.500 -4.000 405.060 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 67.630 -4.000 68.190 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 422.230 -4.000 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 439.960 -4.000 440.520 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 457.690 -4.000 458.250 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 475.420 -4.000 475.980 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 493.150 -4.000 493.710 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 510.880 -4.000 511.440 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 528.610 -4.000 529.170 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 546.340 -4.000 546.900 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 564.070 -4.000 564.630 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 581.800 -4.000 582.360 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 91.270 -4.000 91.830 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 599.530 -4.000 600.090 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 617.260 -4.000 617.820 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 114.910 -4.000 115.470 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 138.550 -4.000 139.110 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 156.280 -4.000 156.840 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 174.010 -4.000 174.570 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 191.740 -4.000 192.300 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 209.470 -4.000 210.030 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 227.200 -4.000 227.760 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 49.900 -4.000 50.460 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 250.840 -4.000 251.400 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 268.570 -4.000 269.130 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 286.300 -4.000 286.860 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 304.030 -4.000 304.590 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 321.760 -4.000 322.320 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 339.490 -4.000 340.050 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 357.220 -4.000 357.780 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 374.950 -4.000 375.510 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 392.680 -4.000 393.240 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 410.410 -4.000 410.970 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 73.540 -4.000 74.100 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 428.140 -4.000 428.700 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 445.870 -4.000 446.430 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 463.600 -4.000 464.160 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 481.330 -4.000 481.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 499.060 -4.000 499.620 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 516.790 -4.000 517.350 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 534.520 -4.000 535.080 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 552.250 -4.000 552.810 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 569.980 -4.000 570.540 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 587.710 -4.000 588.270 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 97.180 -4.000 97.740 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 605.440 -4.000 606.000 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 623.170 -4.000 623.730 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 120.820 -4.000 121.380 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 144.460 -4.000 145.020 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 162.190 -4.000 162.750 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 179.920 -4.000 180.480 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 197.650 -4.000 198.210 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 215.380 -4.000 215.940 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 233.110 -4.000 233.670 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 55.810 -4.000 56.370 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 79.450 -4.000 80.010 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 103.090 -4.000 103.650 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 126.730 -4.000 127.290 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 26.260 -4.000 26.820 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 32.170 -4.000 32.730 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 1728.740 3094.200 1855.470 3145.160 ;
      LAYER met1 ;
        RECT 1730.190 3094.210 1853.575 3147.285 ;
      LAYER met2 ;
        RECT 1730.175 3094.205 1853.590 3147.285 ;
      LAYER met3 ;
        RECT 67.030 3452.485 854.070 3471.460 ;
        RECT 865.870 3452.485 866.570 3471.460 ;
        RECT 878.370 3452.650 1112.570 3471.460 ;
        RECT 1124.370 3452.650 1125.070 3471.460 ;
        RECT 1136.870 3452.650 1594.570 3471.460 ;
        RECT 878.370 3452.485 1594.570 3452.650 ;
        RECT 67.030 3247.050 1594.570 3452.485 ;
        RECT 1620.370 3452.565 1621.070 3471.460 ;
        RECT 1632.870 3460.060 1633.570 3471.460 ;
        RECT 1645.370 3460.060 1646.070 3471.460 ;
        RECT 1632.870 3452.565 1646.070 3460.060 ;
        RECT 1620.370 3247.050 1646.070 3452.565 ;
        RECT 1671.870 3452.400 2552.570 3471.460 ;
        RECT 2577.370 3452.400 2602.570 3471.460 ;
        RECT 2627.370 3452.400 2898.095 3471.460 ;
        RECT 1671.870 3422.080 2898.095 3452.400 ;
        RECT 1671.870 3247.050 2552.570 3422.080 ;
        RECT 67.030 3187.405 2552.570 3247.050 ;
        RECT 2577.370 3223.320 2898.095 3422.080 ;
        RECT 2577.370 3198.520 2833.230 3223.320 ;
        RECT 2577.370 3187.405 2898.095 3198.520 ;
        RECT 67.030 3173.320 2898.095 3187.405 ;
        RECT 67.030 3148.520 2833.230 3173.320 ;
        RECT 67.030 2777.210 2898.095 3148.520 ;
        RECT 67.030 2752.410 2811.195 2777.210 ;
        RECT 67.030 2727.210 2898.095 2752.410 ;
        RECT 67.030 2702.410 2811.195 2727.210 ;
        RECT 67.030 2558.610 2898.095 2702.410 ;
        RECT 1700.760 2557.250 2898.095 2558.610 ;
        RECT 67.030 2501.210 2898.095 2557.250 ;
        RECT 67.030 2499.850 2897.695 2501.210 ;
        RECT 67.030 2495.300 2898.095 2499.850 ;
        RECT 67.030 2493.940 2697.070 2495.300 ;
        RECT 67.030 2318.860 2898.095 2493.940 ;
        RECT 1705.795 2317.500 2898.095 2318.860 ;
        RECT 67.030 2312.950 2898.095 2317.500 ;
        RECT 69.885 2311.590 2898.095 2312.950 ;
        RECT 67.030 2279.100 2898.095 2311.590 ;
        RECT 67.030 2277.740 2897.695 2279.100 ;
        RECT 67.030 2273.190 2898.095 2277.740 ;
        RECT 67.030 2271.830 2686.480 2273.190 ;
        RECT 67.030 2102.750 2898.095 2271.830 ;
        RECT 1709.650 2101.390 2898.095 2102.750 ;
        RECT 67.030 2096.840 2898.095 2101.390 ;
        RECT 69.955 2095.480 2898.095 2096.840 ;
        RECT 67.030 2027.440 2898.095 2095.480 ;
        RECT 67.030 2026.080 2667.085 2027.440 ;
        RECT 67.030 981.550 2898.095 2026.080 ;
        RECT 67.030 957.150 86.705 981.550 ;
        RECT 2868.425 957.150 2882.745 981.550 ;
      LAYER met4 ;
        RECT 69.055 955.490 2884.080 3453.685 ;
      LAYER met5 ;
        RECT 1728.910 2985.260 1854.855 3249.955 ;
  END
END DIGITALTBD
END LIBRARY

